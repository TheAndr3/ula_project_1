module unidade_or_4bits (
    input  wire [3:0] A,    
    input  wire [3:0] B,    
    output wire [3:0] S     
);

    
    or OR0 (S[0], A[0], B[0]);
    or OR1 (S[1], A[1], B[1]);
    or OR2 (S[2], A[2], B[2]);
    or OR3 (S[3], A[3], B[3]);

endmodule
