module mutiplicacao_5x4 (
	input wire [4:0] a,
	input wire [3:0] b,
	output wire [7:0] s

);
	
	wire gnd = 1'b0;
	wire cout01, cout02, cout03, cout04, cout05, cout11, cout12, cout13, cout14, cout15, cout21, cout22, cout23, cout24, cout25;
	wire soma_02;
	//s0
	and U_s0 (s[0], a[0], b[0]);
	
	//s1
	wire b0a1_and, a0b1_and;
	and f0s1 (b0a1_and, a[1], b[0]);
	and f1s1 (a0b1_and, a[0], b[1]);
	
	full_adder soma01 (
	b0a1_and, a0b1_and, gnd,
	s[1], cout01
	);
	
	//s2
	wire a2b0_and, a1b1_and, a0b2_and;

	and f0s2 (a2b0_and, a[2], b[0]);
	and f1s2 (a1b1_and, a[1], b[1]);
	full_adder soma02 (
	a2b0_and, a1b1_and, cout01,
	soma_02, cout02
	);
	and f2s2 (a0b2_and, a[0], b[2]);
	full_adder soma11 (
	a0b2_and, soma_2, gnd,
	s[2], cout11
	);
	
	//s3
	wire a3b0_and, a2b1_and, a1b2_and, a0b3_and;
	wire soma_03, soma_12;
	and f0s3 (a3b0_and, a[3], b[0]);
	and f1s3 (a2b1_and, a[2], b[1]);
	full_adder soma03 (
	a3b0_and, a2b1_and, cout02,
	soma_03, cout03
	);
	and f2s3 (a1b2_and, a[1], b[2]);
	full_adder soma12 (
	a1b2_and, soma_03, cout11,
	soma_12, cout12
	);
	and f3s3 (a0b3_and, a[0], b[3]);
	full_adder soma21 (
	a0b3_and, soma_12, gnd,
	s[3], cout21
	);

	//s4
	wire a4b0_and, a3b1_and, a2b2_and, a1b3_and;
	wire soma_04, soma_13;
	
	and f0s4 (a4b0_and, a[4], b[0]);
	and f1s4 (a3b1_and, a[3], b[1]);
	full_adder soma04 (
	a4b0_and, a3b1_and, cout03,
	soma_04, cout04
	);
	and f2s4 (a2b2_and, a[2], b[2]);
	full_adder soma13 (
	a2b2_and, soma_04, cout12,
	soma_13, cout13
	);
	and f3s4 (a1b3_and, a[1], b[3]);
	full_adder soma22 (
	a1b3_and, soma_13, cout21,
	s[4], cout22
	);
	
	//s5
	wire a4b1_and, a3b2_and, a2b3_and ;
	wire soma_05, soma_14;
	
	and f0s5 (a4b1_and, a[4], b[1]);
	full_adder soma05 (
	a4b1_and, cout04, gnd,
	soma_05, cout05
	);
	and f1s5 (a3b2_and, a[3], b[2]);
	full_adder soma14 (
	a3b2_and, soma_05, cout13,
	soma_14, cout14
	);
	and f2s5 (a2b3_and, a[2], b[3]);
	full_adder soma23 (
	a2b3_and, soma_14, cout22,
	s[5], cout23
	);
	
	//s6
	wire a4b2_and, a3b3_and;
	wire soma_15;
	
	and f0s6 (a4b2_and, a[4], b[2]);
	full_adder soma15 (
	a4b2_and, cout05, cout14,
	soma_15, cout15
	);
	and f1s6 (a3b3_and, a[3], b[3]);
	full_adder soma24 (
	a3b3_and, soma_15, cout23,
	s[6], cout24
	);
	
	//s7
	wire a4b3_and;
	
	and f0s7 (a4b3_and, a[4], b[3]);
	full_adder soma25 (
	a4b3_and, cout15, cout24,
	s[7], cout25
	);


endmodule